(* blackbox *)
module and2(input A1, A2, output Z);
endmodule

(* blackbox *)
module xor2(input A1, A2, output Z);
endmodule

(* blackbox *)
module inv(input I, output ZN);
endmodule

(* blackbox *)
module addf(input A, B, CI, output CO, S);
endmodule

(* blackbox *)
module addh(input A, B, output CO, S);
endmodule

(* blackbox *)
module ao21(input A1, A2, B, output Z);
endmodule

(* blackbox *)
module ao22(input A1, A2, B1, B2, output Z);
endmodule

(* blackbox *)
module oai33(input A1, A2, A3, B1, B2, B3, output ZN);
endmodule
